// This version replaces the enable signal en with a load signal ld. 
// When ld is asserted, the value v is loaded into the counter as a pre-set value.
module counter #(
  parameter WIDTH = 8
)(
  // interface signals
  input  logic             clk,      // clock
  input  logic             rst,      // reset
  input  logic             ld,       // load counter from data
  input  logic [WIDTH-1:0] v,        // value to preload
  output logic [WIDTH-1:0] count     // count output
);

always_ff @ (posedge clk) begin
  if (rst)      count <= {WIDTH{1'b0}};
  else if (ld)  count <= count + 1'b1;
end
endmodule
